

//Model to OR Gate level direct inbuilt function implementation

module orgate_level(output y,input a, inputb);

//input x,y;
//output z;

or(y,a,b);

endmodule