
//Model to OR Gate

module orgate(x,y,z);

input x,y;
output z;

assign z=(x|y);

endmodule
