
//Name: Nuthi Sriram 
//regno: CSE18083

module aluOperations_tb;
reg A,B;
reg [2:0]S;
wire F;
aluOperations dut(.S(S),.A(A),.B(B),.F(F));
initial
 begin
 A=1'b0;
 B=1'b1;
 S=3'b011;
#10
 A=1'b0;
 B=1'b1;
 S=3'b101;
#10
 A=1'b0;
 B=1'b1;
 S=3'b000;
#10
 A=1'b0;
 B=1'b1;
 S=3'b001;
#10
 A=1'b0;
 B=1'b1;
 S=3'b010;
#10
 A=1'b0;
 B=1'b1;
 S=3'b100;
#10
 A=1'b0;
 B=1'b1;
 S=3'b110;
#10
 A=1'b0;
 B=1'b1;
 S=3'b111;
#10
$finish;
end
initial
 $monitor("At time %t, A=%d  B=%d S=%d  =F=%d ", $time,A,B,S,F);
endmodule