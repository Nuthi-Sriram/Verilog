//Implementing a four is to one mux using conditional statements

module fouristoOneMuxUsingConditionalStatement(
input i0, input i1, input i2, input i3, input s0, input s1, output out
);

assign out=s1 ? (s0?i3:i2) : (s0?i1:i0);

endmodule